// QSys.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module QSys (
		input  wire        clk_clk,                    //                 clk.clk
		output wire [10:0] display_buffer_addr_export, // display_buffer_addr.export
		output wire [7:0]  display_buffer_ctrl_export, // display_buffer_ctrl.export
		output wire [31:0] display_buffer_data_export, // display_buffer_data.export
		output wire        epcs_dclk,                  //                epcs.dclk
		output wire        epcs_sce,                   //                    .sce
		output wire        epcs_sdo,                   //                    .sdo
		input  wire        epcs_data0,                 //                    .data0
		output wire [7:0]  pio_led_export,             //             pio_led.export
		input  wire        pll_areset_export,          //          pll_areset.export
		output wire        pll_locked_export,          //          pll_locked.export
		input  wire        reset_reset_n,              //               reset.reset_n
		output wire [12:0] sdram_addr,                 //               sdram.addr
		output wire [1:0]  sdram_ba,                   //                    .ba
		output wire        sdram_cas_n,                //                    .cas_n
		output wire        sdram_cke,                  //                    .cke
		output wire        sdram_cs_n,                 //                    .cs_n
		inout  wire [15:0] sdram_dq,                   //                    .dq
		output wire [1:0]  sdram_dqm,                  //                    .dqm
		output wire        sdram_ras_n,                //                    .ras_n
		output wire        sdram_we_n,                 //                    .we_n
		output wire        sdram_clk_clk,              //           sdram_clk.clk
		output wire        sys_clk_clk,                //             sys_clk.clk
		input  wire        uart_0_rxd,                 //              uart_0.rxd
		output wire        uart_0_txd                  //                    .txd
	);

	wire         cpu_debug_reset_request_reset;                                        // cpu:debug_reset_request -> [display_buffer_addr:reset_n, display_buffer_ctrl:reset_n, display_buffer_data:reset_n, mm_interconnect_0:display_buffer_addr_reset_reset_bridge_in_reset_reset, rst_controller_001:reset_in1, timer_0:reset_n, uart_0:reset_n]
	wire  [31:0] cpu_data_master_readdata;                                             // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                          // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                          // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                              // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                           // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                 // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                                // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                            // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                      // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                   // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                       // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                          // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;               // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;            // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                       // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                        // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                       // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                    // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                    // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                        // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                           // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                     // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                          // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                      // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_controller_epcs_control_port_chipselect -> epcs_flash_controller:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata;   // epcs_flash_controller:readdata -> mm_interconnect_0:epcs_flash_controller_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_controller_epcs_control_port_address -> epcs_flash_controller:address
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_controller_epcs_control_port_read -> epcs_flash_controller:read_n
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_controller_epcs_control_port_write -> epcs_flash_controller:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_controller_epcs_control_port_writedata -> epcs_flash_controller:writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                        // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                         // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                            // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                           // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                       // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                       // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_readdata;                         // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_s1_address;                          // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [1:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                       // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                            // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_writedata;                        // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                            // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_pio_led_s1_chipselect;                              // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                                // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                                 // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                                   // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                               // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;                     // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_readdata;                       // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;                    // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_controller_s1_address;                        // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                           // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controller_s1_byteenable;                     // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;                  // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;                          // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_writedata;                      // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                        // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                          // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                           // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                             // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                         // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_display_buffer_addr_s1_chipselect;                  // mm_interconnect_0:display_buffer_addr_s1_chipselect -> display_buffer_addr:chipselect
	wire  [31:0] mm_interconnect_0_display_buffer_addr_s1_readdata;                    // display_buffer_addr:readdata -> mm_interconnect_0:display_buffer_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_display_buffer_addr_s1_address;                     // mm_interconnect_0:display_buffer_addr_s1_address -> display_buffer_addr:address
	wire         mm_interconnect_0_display_buffer_addr_s1_write;                       // mm_interconnect_0:display_buffer_addr_s1_write -> display_buffer_addr:write_n
	wire  [31:0] mm_interconnect_0_display_buffer_addr_s1_writedata;                   // mm_interconnect_0:display_buffer_addr_s1_writedata -> display_buffer_addr:writedata
	wire         mm_interconnect_0_display_buffer_data_s1_chipselect;                  // mm_interconnect_0:display_buffer_data_s1_chipselect -> display_buffer_data:chipselect
	wire  [31:0] mm_interconnect_0_display_buffer_data_s1_readdata;                    // display_buffer_data:readdata -> mm_interconnect_0:display_buffer_data_s1_readdata
	wire   [1:0] mm_interconnect_0_display_buffer_data_s1_address;                     // mm_interconnect_0:display_buffer_data_s1_address -> display_buffer_data:address
	wire         mm_interconnect_0_display_buffer_data_s1_write;                       // mm_interconnect_0:display_buffer_data_s1_write -> display_buffer_data:write_n
	wire  [31:0] mm_interconnect_0_display_buffer_data_s1_writedata;                   // mm_interconnect_0:display_buffer_data_s1_writedata -> display_buffer_data:writedata
	wire         mm_interconnect_0_display_buffer_ctrl_s1_chipselect;                  // mm_interconnect_0:display_buffer_ctrl_s1_chipselect -> display_buffer_ctrl:chipselect
	wire  [31:0] mm_interconnect_0_display_buffer_ctrl_s1_readdata;                    // display_buffer_ctrl:readdata -> mm_interconnect_0:display_buffer_ctrl_s1_readdata
	wire   [1:0] mm_interconnect_0_display_buffer_ctrl_s1_address;                     // mm_interconnect_0:display_buffer_ctrl_s1_address -> display_buffer_ctrl:address
	wire         mm_interconnect_0_display_buffer_ctrl_s1_write;                       // mm_interconnect_0:display_buffer_ctrl_s1_write -> display_buffer_ctrl:write_n
	wire  [31:0] mm_interconnect_0_display_buffer_ctrl_s1_writedata;                   // mm_interconnect_0:display_buffer_ctrl_s1_writedata -> display_buffer_ctrl:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                              // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                 // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                   // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                               // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                               // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                 // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                  // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                     // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                            // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                    // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                                // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         irq_mapper_receiver0_irq;                                             // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                             // sys_clk_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                             // epcs_flash_controller:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                             // timer_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                             // uart_0:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                                          // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [cpu:reset_n, epcs_flash_controller:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, pio_led:reset_n, rst_translator:in_reset, sdram_controller:reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                               // rst_controller_001:reset_req -> [cpu:reset_req, epcs_flash_controller:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]

	QSys_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_clk_clk),                                  //                    c0.clk
		.c1                 (sys_clk_clk),                                    //                    c1.clk
		.areset             (pll_areset_export),                              //        areset_conduit.export
		.locked             (pll_locked_export),                              //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0),                                           //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0)                                            //           (terminated)
	);

	QSys_cpu cpu (
		.clk                                 (sys_clk_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	QSys_display_buffer_addr display_buffer_addr (
		.clk        (sys_clk_clk),                                         //                 clk.clk
		.reset_n    (~cpu_debug_reset_request_reset),                      //               reset.reset_n
		.address    (mm_interconnect_0_display_buffer_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display_buffer_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display_buffer_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display_buffer_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display_buffer_addr_s1_readdata),   //                    .readdata
		.out_port   (display_buffer_addr_export)                           // external_connection.export
	);

	QSys_display_buffer_ctrl display_buffer_ctrl (
		.clk        (sys_clk_clk),                                         //                 clk.clk
		.reset_n    (~cpu_debug_reset_request_reset),                      //               reset.reset_n
		.address    (mm_interconnect_0_display_buffer_ctrl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display_buffer_ctrl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display_buffer_ctrl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display_buffer_ctrl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display_buffer_ctrl_s1_readdata),   //                    .readdata
		.out_port   (display_buffer_ctrl_export)                           // external_connection.export
	);

	QSys_display_buffer_data display_buffer_data (
		.clk        (sys_clk_clk),                                         //                 clk.clk
		.reset_n    (~cpu_debug_reset_request_reset),                      //               reset.reset_n
		.address    (mm_interconnect_0_display_buffer_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display_buffer_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display_buffer_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display_buffer_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display_buffer_data_s1_readdata),   //                    .readdata
		.out_port   (display_buffer_data_export)                           // external_connection.export
	);

	QSys_epcs_flash_controller epcs_flash_controller (
		.clk        (sys_clk_clk),                                                          //               clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                                  //             reset.reset_n
		.reset_req  (rst_controller_001_reset_out_reset_req),                               //                  .reset_req
		.address    (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver2_irq),                                             //               irq.irq
		.dclk       (epcs_dclk),                                                            //          external.export
		.sce        (epcs_sce),                                                             //                  .export
		.sdo        (epcs_sdo),                                                             //                  .export
		.data0      (epcs_data0)                                                            //                  .export
	);

	QSys_jtag_uart jtag_uart (
		.clk            (sys_clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	QSys_onchip_memory2 onchip_memory2 (
		.clk        (sys_clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	QSys_display_buffer_ctrl pio_led (
		.clk        (sys_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_export)                           // external_connection.export
	);

	QSys_sdram_controller sdram_controller (
		.clk            (sys_clk_clk),                                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	QSys_sys_clk_timer sys_clk_timer (
		.clk        (sys_clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                       //   irq.irq
	);

	QSys_sysid sysid (
		.clock    (sys_clk_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	QSys_sys_clk_timer timer_0 (
		.clk        (sys_clk_clk),                             //   clk.clk
		.reset_n    (~cpu_debug_reset_request_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	QSys_uart_0 uart_0 (
		.clk           (sys_clk_clk),                               //                 clk.clk
		.reset_n       (~cpu_debug_reset_request_reset),            //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_rxd),                                // external_connection.export
		.txd           (uart_0_txd),                                //                    .export
		.irq           (irq_mapper_receiver4_irq)                   //                 irq.irq
	);

	QSys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c1_clk                                            (sys_clk_clk),                                                          //                                          altpll_0_c1.clk
		.clk_50_clk_clk                                             (clk_clk),                                                              //                                           clk_50_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                       // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),                                   //                      cpu_reset_reset_bridge_in_reset.reset
		.display_buffer_addr_reset_reset_bridge_in_reset_reset      (cpu_debug_reset_request_reset),                                        //      display_buffer_addr_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                    (cpu_data_master_address),                                              //                                      cpu_data_master.address
		.cpu_data_master_waitrequest                                (cpu_data_master_waitrequest),                                          //                                                     .waitrequest
		.cpu_data_master_byteenable                                 (cpu_data_master_byteenable),                                           //                                                     .byteenable
		.cpu_data_master_read                                       (cpu_data_master_read),                                                 //                                                     .read
		.cpu_data_master_readdata                                   (cpu_data_master_readdata),                                             //                                                     .readdata
		.cpu_data_master_write                                      (cpu_data_master_write),                                                //                                                     .write
		.cpu_data_master_writedata                                  (cpu_data_master_writedata),                                            //                                                     .writedata
		.cpu_data_master_debugaccess                                (cpu_data_master_debugaccess),                                          //                                                     .debugaccess
		.cpu_instruction_master_address                             (cpu_instruction_master_address),                                       //                               cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                         (cpu_instruction_master_waitrequest),                                   //                                                     .waitrequest
		.cpu_instruction_master_read                                (cpu_instruction_master_read),                                          //                                                     .read
		.cpu_instruction_master_readdata                            (cpu_instruction_master_readdata),                                      //                                                     .readdata
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                         //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                           //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                            //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                        //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                       //                                                     .writedata
		.cpu_debug_mem_slave_address                                (mm_interconnect_0_cpu_debug_mem_slave_address),                        //                                  cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                  (mm_interconnect_0_cpu_debug_mem_slave_write),                          //                                                     .write
		.cpu_debug_mem_slave_read                                   (mm_interconnect_0_cpu_debug_mem_slave_read),                           //                                                     .read
		.cpu_debug_mem_slave_readdata                               (mm_interconnect_0_cpu_debug_mem_slave_readdata),                       //                                                     .readdata
		.cpu_debug_mem_slave_writedata                              (mm_interconnect_0_cpu_debug_mem_slave_writedata),                      //                                                     .writedata
		.cpu_debug_mem_slave_byteenable                             (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                     //                                                     .byteenable
		.cpu_debug_mem_slave_waitrequest                            (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                    //                                                     .waitrequest
		.cpu_debug_mem_slave_debugaccess                            (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                    //                                                     .debugaccess
		.display_buffer_addr_s1_address                             (mm_interconnect_0_display_buffer_addr_s1_address),                     //                               display_buffer_addr_s1.address
		.display_buffer_addr_s1_write                               (mm_interconnect_0_display_buffer_addr_s1_write),                       //                                                     .write
		.display_buffer_addr_s1_readdata                            (mm_interconnect_0_display_buffer_addr_s1_readdata),                    //                                                     .readdata
		.display_buffer_addr_s1_writedata                           (mm_interconnect_0_display_buffer_addr_s1_writedata),                   //                                                     .writedata
		.display_buffer_addr_s1_chipselect                          (mm_interconnect_0_display_buffer_addr_s1_chipselect),                  //                                                     .chipselect
		.display_buffer_ctrl_s1_address                             (mm_interconnect_0_display_buffer_ctrl_s1_address),                     //                               display_buffer_ctrl_s1.address
		.display_buffer_ctrl_s1_write                               (mm_interconnect_0_display_buffer_ctrl_s1_write),                       //                                                     .write
		.display_buffer_ctrl_s1_readdata                            (mm_interconnect_0_display_buffer_ctrl_s1_readdata),                    //                                                     .readdata
		.display_buffer_ctrl_s1_writedata                           (mm_interconnect_0_display_buffer_ctrl_s1_writedata),                   //                                                     .writedata
		.display_buffer_ctrl_s1_chipselect                          (mm_interconnect_0_display_buffer_ctrl_s1_chipselect),                  //                                                     .chipselect
		.display_buffer_data_s1_address                             (mm_interconnect_0_display_buffer_data_s1_address),                     //                               display_buffer_data_s1.address
		.display_buffer_data_s1_write                               (mm_interconnect_0_display_buffer_data_s1_write),                       //                                                     .write
		.display_buffer_data_s1_readdata                            (mm_interconnect_0_display_buffer_data_s1_readdata),                    //                                                     .readdata
		.display_buffer_data_s1_writedata                           (mm_interconnect_0_display_buffer_data_s1_writedata),                   //                                                     .writedata
		.display_buffer_data_s1_chipselect                          (mm_interconnect_0_display_buffer_data_s1_chipselect),                  //                                                     .chipselect
		.epcs_flash_controller_epcs_control_port_address            (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    //              epcs_flash_controller_epcs_control_port.address
		.epcs_flash_controller_epcs_control_port_write              (mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),      //                                                     .write
		.epcs_flash_controller_epcs_control_port_read               (mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),       //                                                     .read
		.epcs_flash_controller_epcs_control_port_readdata           (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                                                     .readdata
		.epcs_flash_controller_epcs_control_port_writedata          (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                                                     .writedata
		.epcs_flash_controller_epcs_control_port_chipselect         (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                                                     .chipselect
		.jtag_uart_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                //                          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                  //                                                     .write
		.jtag_uart_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                   //                                                     .read
		.jtag_uart_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),               //                                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),              //                                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),            //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),             //                                                     .chipselect
		.onchip_memory2_s1_address                                  (mm_interconnect_0_onchip_memory2_s1_address),                          //                                    onchip_memory2_s1.address
		.onchip_memory2_s1_write                                    (mm_interconnect_0_onchip_memory2_s1_write),                            //                                                     .write
		.onchip_memory2_s1_readdata                                 (mm_interconnect_0_onchip_memory2_s1_readdata),                         //                                                     .readdata
		.onchip_memory2_s1_writedata                                (mm_interconnect_0_onchip_memory2_s1_writedata),                        //                                                     .writedata
		.onchip_memory2_s1_byteenable                               (mm_interconnect_0_onchip_memory2_s1_byteenable),                       //                                                     .byteenable
		.onchip_memory2_s1_chipselect                               (mm_interconnect_0_onchip_memory2_s1_chipselect),                       //                                                     .chipselect
		.onchip_memory2_s1_clken                                    (mm_interconnect_0_onchip_memory2_s1_clken),                            //                                                     .clken
		.pio_led_s1_address                                         (mm_interconnect_0_pio_led_s1_address),                                 //                                           pio_led_s1.address
		.pio_led_s1_write                                           (mm_interconnect_0_pio_led_s1_write),                                   //                                                     .write
		.pio_led_s1_readdata                                        (mm_interconnect_0_pio_led_s1_readdata),                                //                                                     .readdata
		.pio_led_s1_writedata                                       (mm_interconnect_0_pio_led_s1_writedata),                               //                                                     .writedata
		.pio_led_s1_chipselect                                      (mm_interconnect_0_pio_led_s1_chipselect),                              //                                                     .chipselect
		.sdram_controller_s1_address                                (mm_interconnect_0_sdram_controller_s1_address),                        //                                  sdram_controller_s1.address
		.sdram_controller_s1_write                                  (mm_interconnect_0_sdram_controller_s1_write),                          //                                                     .write
		.sdram_controller_s1_read                                   (mm_interconnect_0_sdram_controller_s1_read),                           //                                                     .read
		.sdram_controller_s1_readdata                               (mm_interconnect_0_sdram_controller_s1_readdata),                       //                                                     .readdata
		.sdram_controller_s1_writedata                              (mm_interconnect_0_sdram_controller_s1_writedata),                      //                                                     .writedata
		.sdram_controller_s1_byteenable                             (mm_interconnect_0_sdram_controller_s1_byteenable),                     //                                                     .byteenable
		.sdram_controller_s1_readdatavalid                          (mm_interconnect_0_sdram_controller_s1_readdatavalid),                  //                                                     .readdatavalid
		.sdram_controller_s1_waitrequest                            (mm_interconnect_0_sdram_controller_s1_waitrequest),                    //                                                     .waitrequest
		.sdram_controller_s1_chipselect                             (mm_interconnect_0_sdram_controller_s1_chipselect),                     //                                                     .chipselect
		.sys_clk_timer_s1_address                                   (mm_interconnect_0_sys_clk_timer_s1_address),                           //                                     sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                                     (mm_interconnect_0_sys_clk_timer_s1_write),                             //                                                     .write
		.sys_clk_timer_s1_readdata                                  (mm_interconnect_0_sys_clk_timer_s1_readdata),                          //                                                     .readdata
		.sys_clk_timer_s1_writedata                                 (mm_interconnect_0_sys_clk_timer_s1_writedata),                         //                                                     .writedata
		.sys_clk_timer_s1_chipselect                                (mm_interconnect_0_sys_clk_timer_s1_chipselect),                        //                                                     .chipselect
		.sysid_control_slave_address                                (mm_interconnect_0_sysid_control_slave_address),                        //                                  sysid_control_slave.address
		.sysid_control_slave_readdata                               (mm_interconnect_0_sysid_control_slave_readdata),                       //                                                     .readdata
		.timer_0_s1_address                                         (mm_interconnect_0_timer_0_s1_address),                                 //                                           timer_0_s1.address
		.timer_0_s1_write                                           (mm_interconnect_0_timer_0_s1_write),                                   //                                                     .write
		.timer_0_s1_readdata                                        (mm_interconnect_0_timer_0_s1_readdata),                                //                                                     .readdata
		.timer_0_s1_writedata                                       (mm_interconnect_0_timer_0_s1_writedata),                               //                                                     .writedata
		.timer_0_s1_chipselect                                      (mm_interconnect_0_timer_0_s1_chipselect),                              //                                                     .chipselect
		.uart_0_s1_address                                          (mm_interconnect_0_uart_0_s1_address),                                  //                                            uart_0_s1.address
		.uart_0_s1_write                                            (mm_interconnect_0_uart_0_s1_write),                                    //                                                     .write
		.uart_0_s1_read                                             (mm_interconnect_0_uart_0_s1_read),                                     //                                                     .read
		.uart_0_s1_readdata                                         (mm_interconnect_0_uart_0_s1_readdata),                                 //                                                     .readdata
		.uart_0_s1_writedata                                        (mm_interconnect_0_uart_0_s1_writedata),                                //                                                     .writedata
		.uart_0_s1_begintransfer                                    (mm_interconnect_0_uart_0_s1_begintransfer),                            //                                                     .begintransfer
		.uart_0_s1_chipselect                                       (mm_interconnect_0_uart_0_s1_chipselect)                                //                                                     .chipselect
	);

	QSys_irq_mapper irq_mapper (
		.clk           (sys_clk_clk),                        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.clk            (sys_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
